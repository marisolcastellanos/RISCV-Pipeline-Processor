module if_id( 
              input logic clk,reset, 
              input 
