module idecode ( 
                input  logic        clk,reset,
                input  logic [31:0] InstrD, 
                input  logic [31:0] PCD, PCPlus4D,
                input  logic        RegWriteW,
                input  logic        ResultW,
                input  logic        RdW,
                );
endmodule
